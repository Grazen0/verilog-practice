`ifndef _NOTES_VH_
`define _NOTES_VH_

`define NOTE(note, duration) ((((duration) & 4'hF) << 8) | ((note) & 8'hFF))
`define TO_DIVIDER(clk, freq) (clk) / (2 * (freq))

`define SILENCE 0
`define C0 1
`define CS0 2
`define D0 3
`define EB0 4
`define E0 5
`define F0 6
`define FS0 7
`define G0 8
`define AB0 9
`define A0 10
`define BB0 11
`define B0 12
`define C1 13
`define CS1 14
`define D1 15
`define EB1 16
`define E1 17
`define F1 18
`define FS1 19
`define G1 20
`define AB1 21
`define A1 22
`define BB1 23
`define B1 24
`define C2 25
`define CS2 26
`define D2 27
`define EB2 28
`define E2 29
`define F2 30
`define FS2 31
`define G2 32
`define AB2 33
`define A2 34
`define BB2 35
`define B2 36
`define C3 37
`define CS3 38
`define D3 39
`define EB3 40
`define E3 41
`define F3 42
`define FS3 43
`define G3 44
`define AB3 45
`define A3 46
`define BB3 47
`define B3 48
`define C4 49
`define CS4 50
`define D4 51
`define EB4 52
`define E4 53
`define F4 54
`define FS4 55
`define G4 56
`define AB4 57
`define A4 58
`define BB4 59
`define B4 60
`define C5 61
`define CS5 62
`define D5 63
`define EB5 64
`define E5 65
`define F5 66
`define FS5 67
`define G5 68
`define AB5 69
`define A5 70
`define BB5 71
`define B5 72
`define C6 73
`define CS6 74
`define D6 75
`define EB6 76
`define E6 77
`define F6 78
`define FS6 79
`define G6 80
`define AB6 81
`define A6 82
`define BB6 83
`define B6 84
`define C7 85
`define CS7 86
`define D7 87
`define EB7 88
`define E7 89
`define F7 90
`define FS7 91
`define G7 92
`define AB7 93
`define A7 94
`define BB7 95
`define B7 96
`define C8 97
`define CS8 98
`define D8 99
`define EB8 100
`define E8 101
`define F8 102
`define FS8 103
`define G8 104
`define AB8 105
`define A8 106
`define BB8 107
`define B8 108

`endif
