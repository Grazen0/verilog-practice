module music_player ();

endmodule
